//package ibex_dv_pkg;
        `include "dv_macros.svh"
	`include "bus_params_pkg.sv"
	`include "common_ifs_pkg.sv"
	`include "clk_rst_if.sv"
	`include "irq_if.sv"
	`include "ibex_mem_intf.sv"
	`include "str_utils_pkg.sv"
	`include "dv_utils_pkg.sv"
       	`include "../rtl/ibex_pkg.sv"
	`include "core_ibex_dut_probe_if.sv"
	`include "core_ibex_instr_monitor_if.sv"
	`include "core_ibex_rvfi_if.sv"
	`include "core_ibex_csr_if.sv"
	`include "core_ibex_ifetch_if.sv"
	`include "core_ibex_ifetch_pmp_if.sv"
	`include "push_pull_if.sv"
	//`include "prim_secded_pkg.sv"
	//`include "irq_agent_pkg.sv"
	`include "ibex_mem_intf_pkg.sv"
	//`include "ibex_cosim_agent_pkg.sv"
//endpackage
